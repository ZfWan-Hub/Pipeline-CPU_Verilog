`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:45:02 11/16/2018 
// Design Name: 
// Module Name:    DM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DM(
    input [9:0] Addr,
    input [31:0] DataIn,
    input DMwrite,
	 input [31:0]PC,
    input clk,
    input reset,
    output [31:0] DataOut
    );

	reg [31:0] dm_reg [1023:0];
	integer i;
	
	initial begin
		for(i=0;i<1024;i=i+1)begin
				dm_reg[i]=0;
			end
	end
	
	assign DataOut= dm_reg[Addr];
	
	always@(posedge clk )begin
		if(reset)begin
			for(i=0;i<1024;i=i+1)begin
				dm_reg[i]=0;
			end
		end
		else begin
			if(DMwrite)begin
				dm_reg[Addr]=DataIn;
				$display("@%h: *%h <= %h",PC, {20'd0,Addr,2'b0},DataIn); 
			end
		end
	end
endmodule
